player entities/columbiare 803 150
world world/world.wld
npc stand entities/npcs/test.npc
npc stand entities/npcs/amia.npc
npc stand entities/npcs/fara.npc
progress a1s1